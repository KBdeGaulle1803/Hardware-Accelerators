`timescale 1ns / 1ps

module PLAN_ctrl(
input [31:0] num,
input clk, res,
output reg [31:0] x, cf1, cf2
);
reg posres;

always@(posedge clk)
begin
x=(res)?32'd0:num;

if(res) cf1=32'd0;
else if(x[30:23]<8'd125) cf1=(x[31])?32'h3E7ECE00:32'hBE7ECE00;
else if(x[30:23]==8'd125) cf1=(x[31])?32'h3E770A00:32'hBE770A00;
else if(x[30:22]=={8'd126,1'b0}) cf1=(x[31])?32'h3E686E00:32'hBE686E00;
else if(x[30:22]=={8'd126,1'b1}) cf1=(x[31])?32'h3E548700:32'hBE548700;
else if(x[30:21]=={8'd127,2'b00}) cf1=(x[31])?32'h3E3D6C00:32'hBE3D6C00;
else if(x[30:21]=={8'd127,2'b01}) cf1=(x[31])?32'h3E250600:32'hBE250600;
else if(x[30:21]=={8'd127,2'b10}) cf1=(x[31])?32'h3E0CC500:32'hBE0CC500;
else if(x[30:21]=={8'd127,2'b11}) cf1=(x[31])?32'h3DEC5000:32'hBDEC5000;
else if(x[30:20]=={8'd128,3'b000}) cf1=(x[31])?32'h3DC35000:32'hBDC35000;
else if(x[30:20]=={8'd128,3'b001}) cf1=(x[31])?32'h3D9F9000:32'hBD9F9000;
else if(x[30:20]=={8'd128,3'b010}) cf1=(x[31])?32'h3D812200:32'hBD812200;
else if(x[30:20]=={8'd128,3'b011}) cf1=(x[31])?32'h3D4F5000:32'hBD4F5000;
else if(x[30:20]=={8'd128,3'b100}) cf1=(x[31])?32'h3D254000:32'hBD254000;
else if(x[30:20]=={8'd128,3'b101}) cf1=(x[31])?32'h3D033000:32'hBD033000;
else if(x[30:20]=={8'd128,3'b110}) cf1=(x[31])?32'h3CCF8000:32'hBCCF8000;
else if(x[30:20]=={8'd128,3'b111}) cf1=(x[31])?32'h3CA35800:32'hBCA35800;
else if(x[30:19]=={8'd129,4'b0000}) cf1=(x[31])?32'h3C805E00:32'hBC805E00;
else if(x[30:19]=={8'd129,4'b0001}) cf1=(x[31])?32'h3C497400:32'hBC497400;
else if(x[30:19]=={8'd129,4'b0010}) cf1=(x[31])?32'h3C1DB400:32'hBC1DB400;
else if(x[30:19]=={8'd129,4'b0011}) cf1=(x[31])?32'h3BF6FC00:32'hBBF6FC00;
else if(x[30:19]=={8'd129,4'b0100}) cf1=(x[31])?32'h3BC0CC00:32'hBBC0CC00;
else if(x[30:19]=={8'd129,4'b0101}) cf1=(x[31])?32'h3B968400:32'hBB968400;
else if(x[30:19]=={8'd129,4'b0110}) cf1=(x[31])?32'h3B6AC000:32'hBB6AC000;
else if(x[30:19]=={8'd129,4'b0111}) cf1=(x[31])?32'h3B373800:32'hBB373800;
else if(x[30:19]=={8'd129,4'b1000}) cf1=(x[31])?32'h3B0EE400:32'hBB0EE400;
else if(x[30:19]=={8'd129,4'b1001}) cf1=(x[31])?32'h3ADDC931:32'hBADDC931;
else if(x[30:19]=={8'd129,4'b1010}) cf1=(x[31])?32'h3AAD8000:32'hBAAD8000;
else if(x[30:19]=={8'd129,4'b1011}) cf1=(x[31])?32'h3A876400:32'hBA876400;
else if(x[30:19]=={8'd129,4'b1100}) cf1=(x[31])?32'h3A52E800:32'hBA52E800;
else if(x[30:19]=={8'd129,4'b1101}) cf1=(x[31])?32'h3A24AC03:32'hBA24AC03;
else if(x[30:19]=={8'd129,4'b1110}) cf1=(x[31])?32'h39FF9800:32'hB9FF9800;
else if(x[30:19]=={8'd129,4'b1111}) cf1=(x[31])?32'h39C76800:32'hB9C76800;
else if(x[30:18]=={8'd130,5'b00000}) cf1=(x[31])?32'h399BC800:32'hB99BC800;
else if(x[30:18]=={8'd130,5'b00001}) cf1=(x[31])?32'h39723000:32'hB9723000;
else if(x[30:18]=={8'd130,5'b00010}) cf1=(x[31])?32'h393CE000:32'hB93CE000;
else if(x[30:18]=={8'd130,5'b00011}) cf1=(x[31])?32'h3912F400:32'hB912F400;
else if(x[30:18]=={8'd130,5'b00100}) cf1=(x[31])?32'h38E52800:32'hB8E52800;
else if(x[30:18]=={8'd130,5'b00101}) cf1=(x[31])?32'h38B267FF:32'hB8B267FF;
else if(x[30:18]=={8'd130,5'b00110}) cf1=(x[31])?32'h388AE000:32'hB88AE000;
else if(x[30:18]=={8'd130,5'b00111}) cf1=(x[31])?32'h385BC000:32'hB85BC000;
else if(x[30:18]=={8'd130,5'b01000}) cf1=(x[31])?32'h3828D801:32'hB828D801;
else if(x[30:18]=={8'd130,5'b01001}) cf1=(x[31])?32'h38033000:32'hB8033000;
else if(x[30:18]=={8'd130,5'b01010}) cf1=(x[31])?32'h37CC67FF:32'hB7CC67FF;
else if(x[30:18]=={8'd130,5'b01011}) cf1=(x[31])?32'h379F4800:32'hB79F4800;
else if(x[30:18]=={8'd130,5'b01100}) cf1=(x[31])?32'h37783000:32'hB7783000;
else if(x[30:18]=={8'd130,5'b01101}) cf1=(x[31])?32'h3740D801:32'hB740D801;
else if(x[30:18]=={8'd130,5'b01110}) cf1=(x[31])?32'h37169000:32'hB7169000;
else if(x[30:18]=={8'd130,5'b01111}) cf1=(x[31])?32'h36EB3000:32'hB6EB3000;
else if(x[30:18]=={8'd130,5'b10000}) cf1=(x[31])?32'h36B67000:32'hB6B67000;
else if(x[30:18]=={8'd130,5'b10001}) cf1=(x[31])?32'h368D9000:32'hB68D9000;
else if(x[30:18]=={8'd130,5'b10010}) cf1=(x[31])?32'h365DE001:32'hB65DE001;
else if(x[30:18]=={8'd130,5'b10011}) cf1=(x[31])?32'h362C6001:32'hB62C6001;
else if(x[30:18]=={8'd130,5'b10100}) cf1=(x[31])?32'h3605B000:32'hB605B000;
else if(x[30:18]=={8'd130,5'b10101}) cf1=(x[31])?32'h35D2D687:32'hB5D2D687;
else if(x[30:18]=={8'd130,5'b10110}) cf1=(x[31])?32'h35A2C000:32'hB5A2C000;
else if(x[30:18]=={8'd130,5'b10111}) cf1=(x[31])?32'h357FD000:32'hB57FD000;
else if(x[30:18]=={8'd130,5'b11000}) cf1=(x[31])?32'h3545E000:32'hB545E000;
else if(x[30:18]=={8'd130,5'b11001}) cf1=(x[31])?32'h351A3000:32'hB51A3000;
else if(x[30:18]=={8'd130,5'b11010}) cf1=(x[31])?32'h34F07000:32'hB4F07000;
else if(x[30:18]=={8'd130,5'b11011}) cf1=(x[31])?32'h34BB3000:32'hB4BB3000;
else if(x[30:18]=={8'd130,5'b11100}) cf1=(x[31])?32'h34923800:32'hB4923800;
else if(x[30:18]=={8'd130,5'b11101}) cf1=(x[31])?32'h34622000:32'hB4622000;
else if(x[30:18]=={8'd130,5'b11110}) cf1=(x[31])?32'h34308000:32'hB4308000;
else if(x[30:18]=={8'd130,5'b11111}) cf1=(x[31])?32'h34095800:32'hB4095800;
else cf1=(x[31])?32'h00000000:32'h80000000;

posres=res;
end

always@(negedge clk)
begin
if(posres) cf2=32'd0;
else if(x[30:23]<8'd125) cf2=(x[31])?32'h3EFFF77C:32'h3F000442;
else if(x[30:23]==8'd125) cf2=(x[31])?32'h3EFEEF00:32'h3F008880;
else if(x[30:22]=={8'd126,1'b0}) cf2=(x[31])?32'h3EFB3B80:32'h3F026240;
else if(x[30:22]=={8'd126,1'b1}) cf2=(x[31])?32'h3EF3BB00:32'h3F062280;
else if(x[30:21]=={8'd127,2'b00}) cf2=(x[31])?32'h3EE82900:32'h3F0BEB80;
else if(x[30:21]=={8'd127,2'b01}) cf2=(x[31])?32'h3ED8E900:32'h3F138B80;
else if(x[30:21]=={8'd127,2'b10}) cf2=(x[31])?32'h3EC6BB00:32'h3F1CA280;
else if(x[30:21]=={8'd127,2'b11}) cf2=(x[31])?32'h3EB2F600:32'h3F268500;
else if(x[30:20]=={8'd128,3'b000}) cf2=(x[31])?32'h3E9E7C00:32'h3F30C200;
else if(x[30:20]=={8'd128,3'b001}) cf2=(x[31])?32'h3E8A6400:32'h3F3ACE00;
else if(x[30:20]=={8'd128,3'b010}) cf2=(x[31])?32'h3E6ECA00:32'h3F444D80;
else if(x[30:20]=={8'd128,3'b011}) cf2=(x[31])?32'h3E4BD200:32'h3F4D0B80;
else if(x[30:20]=={8'd128,3'b100}) cf2=(x[31])?32'h3E2C5000:32'h3F54EC00;
else if(x[30:20]=={8'd128,3'b101}) cf2=(x[31])?32'h3E10A600:32'h3F5BD680;
else if(x[30:20]=={8'd128,3'b110}) cf2=(x[31])?32'h3DF15400:32'h3F61D580;
else if(x[30:20]=={8'd128,3'b111}) cf2=(x[31])?32'h3DC7FA00:32'h3F6700C0;
else if(x[30:19]=={8'd129,4'b0000}) cf2=(x[31])?32'h3DA50A00:32'h3F6B5EC0;
else if(x[30:19]=={8'd129,4'b0001}) cf2=(x[31])?32'h3D87B200:32'h3F6F09C0;
else if(x[30:19]=={8'd129,4'b0010}) cf2=(x[31])?32'h3D5E3800:32'h3F721C80;
else if(x[30:19]=={8'd129,4'b0011}) cf2=(x[31])?32'h3D359C00:32'h3F74A640;
else if(x[30:19]=={8'd129,4'b0100}) cf2=(x[31])?32'h3D13CA00:32'h3F76C360;
else if(x[30:19]=={8'd129,4'b0101}) cf2=(x[31])?32'h3CF01C00:32'h3F787F20;
else if(x[30:19]=={8'd129,4'b0110}) cf2=(x[31])?32'h3CC29400:32'h3F79EB60;
else if(x[30:19]=={8'd129,4'b0111}) cf2=(x[31])?32'h3C9D8C00:32'h3F7B13A0;
else if(x[30:19]=={8'd129,4'b1000}) cf2=(x[31])?32'h3C7EA400:32'h3F7C0570;
else if(x[30:19]=={8'd129,4'b1001}) cf2=(x[31])?32'h3C4D6800:32'h3F7CCA60;
else if(x[30:19]=={8'd129,4'b1010}) cf2=(x[31])?32'h3C257400:32'h3F7D6A30;
else if(x[30:19]=={8'd129,4'b1011}) cf2=(x[31])?32'h3C054C00:32'h3F7DEAD0;
else if(x[30:19]=={8'd129,4'b1100}) cf2=(x[31])?32'h3BD64400:32'h3F7E5378;
else if(x[30:19]=={8'd129,4'b1101}) cf2=(x[31])?32'h3BAC6400:32'h3F7EA738;
else if(x[30:19]=={8'd129,4'b1110}) cf2=(x[31])?32'h3B89D800:32'h3F7EEC50;
else if(x[30:19]=={8'd129,4'b1111}) cf2=(x[31])?32'h3B5D4000:32'h3F7F22C0;
else if(x[30:18]=={8'd130,5'b00000}) cf2=(x[31])?32'h3B31A800:32'h3F7F4E58;
else if(x[30:18]=={8'd130,5'b00001}) cf2=(x[31])?32'h3B0DEC00:32'h3F7F7214;
else if(x[30:18]=={8'd130,5'b00010}) cf2=(x[31])?32'h3AE33000:32'h3F7F8E68;
else if(x[30:18]=={8'd130,5'b00011}) cf2=(x[31])?32'h3AB56800:32'h3F7FA54C;
else if(x[30:18]=={8'd130,5'b00100}) cf2=(x[31])?32'h3A910000:32'h3F7FB780;
else if(x[30:18]=={8'd130,5'b00101}) cf2=(x[31])?32'h3A676000:32'h3F7FC628;
else if(x[30:18]=={8'd130,5'b00110}) cf2=(x[31])?32'h3A387800:32'h3F7FD1E2;
else if(x[30:18]=={8'd130,5'b00111}) cf2=(x[31])?32'h3A152400:32'h3F7FDAB7;
else if(x[30:18]=={8'd130,5'b01000}) cf2=(x[31])?32'h39EAC800:32'h3F7FE2A7;
else if(x[30:18]=={8'd130,5'b01001}) cf2=(x[31])?32'h39BA8800:32'h3F7FE8AF;
else if(x[30:18]=={8'd130,5'b01010}) cf2=(x[31])?32'h39948800:32'h3F7FED6F;
else if(x[30:18]=={8'd130,5'b01011}) cf2=(x[31])?32'h396C6800:32'h3F7FF13A;
else if(x[30:18]=={8'd130,5'b01100}) cf2=(x[31])?32'h393C1000:32'h3F7FF43F;
else if(x[30:18]=={8'd130,5'b01101}) cf2=(x[31])?32'h39152800:32'h3F7FF6AE;
else if(x[30:18]=={8'd130,5'b01110}) cf2=(x[31])?32'h38EDA000:32'h3F7FF893;
else if(x[30:18]=={8'd130,5'b01111}) cf2=(x[31])?32'h38BD27FF:32'h3F7FFA17;
else if(x[30:18]=={8'd130,5'b10000}) cf2=(x[31])?32'h3895B000:32'h3F7FFB52;
else if(x[30:18]=={8'd130,5'b10001}) cf2=(x[31])?32'h386CC000:32'h3F7FFC4D;
else if(x[30:18]=={8'd130,5'b10010}) cf2=(x[31])?32'h383CE000:32'h3F7FFD0C;
else if(x[30:18]=={8'd130,5'b10011}) cf2=(x[31])?32'h38157800:32'h3F7FFDAA;
else if(x[30:18]=={8'd130,5'b10100}) cf2=(x[31])?32'h37EC2000:32'h3F7FFE28;
else if(x[30:18]=={8'd130,5'b10101}) cf2=(x[31])?32'h37BD4000:32'h3F7FFE86;
else if(x[30:18]=={8'd130,5'b10110}) cf2=(x[31])?32'h3794C800:32'h3F7FFED6;
else if(x[30:18]=={8'd130,5'b10111}) cf2=(x[31])?32'h376DB000:32'h3F7FFF12;
else if(x[30:18]=={8'd130,5'b11000}) cf2=(x[31])?32'h373B0000:32'h3F7FFF45;
else if(x[30:18]=={8'd130,5'b11001}) cf2=(x[31])?32'h37142800:32'h3F7FFF6C;
else if(x[30:18]=={8'd130,5'b11010}) cf2=(x[31])?32'h36EAB001:32'h3F7FFF8B;
else if(x[30:18]=={8'd130,5'b11011}) cf2=(x[31])?32'h36B9B000:32'h3F7FFFA3;
else if(x[30:18]=={8'd130,5'b11100}) cf2=(x[31])?32'h36934800:32'h3F7FFFB6;
else if(x[30:18]=={8'd130,5'b11101}) cf2=(x[31])?32'h36677000:32'h3F7FFFC6;
else if(x[30:18]=={8'd130,5'b11110}) cf2=(x[31])?32'h363757FF:32'h3F7FFFD2;
else if(x[30:18]=={8'd130,5'b11111}) cf2=(x[31])?32'h3610E001:32'h3F7FFFDC;
else cf2=(x[31])?32'h00000000:32'h3F800000;
end

endmodule
